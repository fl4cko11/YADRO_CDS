//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input  [3:0] d0, d1,
  input        sel,
  output [3:0] y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1 (
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);

  // Внутренние сигналы
  logic [3:0] y_temp1;
  logic [3:0] y_temp2;

  // Инстанцирование 2:1 мультиплексоров
  mux_2_1 inst_mux_2_1_helper1 (.d0(d0), .d1(d1), .sel(sel[0]), .y(y_temp1));
  mux_2_1 inst_mux_2_1_helper2 (.d0(d2), .d1(d3), .sel(sel[0]), .y(y_temp2));
  mux_2_1 inst_mux_2_1_main (.d0(y_temp1), .d1(y_temp2), .sel(sel[1]), .y(y));

endmodule
